`define WIDTH 8
//`define trans_number 600	// For coverage
`define trans_number 20
