`define WIDTH 8
`define trans_number 10
