`define WIDTH 8
//`define trans_number 200	// For coverage
`define trans_number 30
