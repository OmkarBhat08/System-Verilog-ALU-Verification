package pkg;
	`include "transaction.sv"
	`include "generator.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "reference_model.sv"
	`include "cscoreboard.sv"
	`include "environment.sv"
	`include "test.sv"
endpackage
