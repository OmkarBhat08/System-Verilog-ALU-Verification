`define WIDTH 8
`define trans_number 1000	// For coverage
//`define trans_number 10
